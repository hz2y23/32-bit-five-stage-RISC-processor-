`define R_Type 				7'b0110011
`define I_Type_Load 		7'b0000011
`define S_Type 				7'b0100011
`define I_Type_calculate 	7'b0010011
`define B_Type 				7'b1100011
`define JAL 				7'b1101111
`define LUI 				7'b0110111