`define EXE_ADD			4'b0000
`define EXE_OR		 	4'b0001
`define EXE_AND		 	4'b0010
`define EXE_XOR		 	4'b0011
`define EXE_SLL		 	4'b0100
`define EXE_SRL		 	4'b0101
`define EXE_SUB		 	4'b0110
`define EXE_SRA		 	4'b0111
`define EXE_SLT		 	4'b1000
`define EXE_LUI		 	4'b1001